module CLA(clk_ram, clk_core, ram_iobus);
	input [31:0] ram_iobus;

endmodule
